Q-1b Open the feedback loop and simulate the opamp

C1 0 3 10n IC=0v  
R1 4 5 10k
R2 5 0 10k
G1 0 3 1 0 10m
E2 4 0 3 0 1
*Giving a step input
Vin 1 0 Pulse(0 1 0 0 30 20 20)
.tran 0.005ms 4ms uic

.control
run
*plotting input and output voltages
plot v(1) v(4)
.endc
.end
