NMOS common source amplifier

.model MN4007 NMOS (Kp=500u Vto=1.5 Lambda=0.01 Gamma=0.6+ Xj=0 Tox=1200n Phi=.6 Rs=0 Rd=0 Cbd=2.0p Cbs=2.0p Pb=.8 Cgso=0.1p Cgdo=0.1p Is=16.64p N=1)

M1 0 1 2 0 MN4007

Vdd 3 0 10v
Vin 1 0 dc 10mv

Rd 3 2 4k
R1 3 1 7.5k
R2 1 0 3.214k

.tran 0.002ms 6ms
.control 
run
plot v(2) v(1)
.endc
.end


