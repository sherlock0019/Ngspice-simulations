Bipolar amplifier

.MODEL Q2N2222A NPN(IS=8.11E-14 BF=205 VAF=113 IKF=0.5 ISE=1.06E-11
+ NE=2 BR=4 VAR=24 IKR=0.225 RB=1.37 RE=0.343 RC=0.137 CJE=2.95E-11
+ TF=3.97E-10 CJC=1.52E-11 TR=8.5E-8 XTB=1.5)

Rc 1 3 5k
R1 1 2 65k
R2 2 0 10k
Re 4 0 2k
VCC 1 0 dc=12
Vin 2 0 dc 0 ac 1 sin(1 0.1 500)
Q1 2 3 4 Q2N2222A
.tran 10u 10m
*.ac dec 10 10 1Meg

.control
run
plot v(2) v(3)
.endc
