Simple voltage regulator circuit using Zener diode
V1 a 0 dc 0 Sin(0 2.5 1k 0 0 0)
Rs a b 1Meg
D1 0 b D1N4148
RL b 0 1Meg

.model D1N4148 D(Is=5.84n N=1.94 Rs=.7017 Ikf=44.17m Xti=3 Eg=1.11 Cjo=.95p M=.55 Vj=.75 Fc=.5 Isr=11.07n Nr=2.088 Bv=100 Ibv=100u Tt=11.07n)
.tran 0.01ms 10ms

*control statements
.control
run

*white background
set color0=white
* black grid and text (only needed with X11, automatic with MS Win)
set color1=black
* wider grid and plot lines
set xbrushwidth=2

plot v(a) v(b)
.endc
.end

