Clipper Circuit

Vin 1 0 DC=0 SIN(0 2.5 1K 0 0)
V1 3 0 dc=2
R1 2 1 1k
D1 2 3 D1N750
*.model D1N750 D(Vj=.75 Cjo=175p Rs=.25 Eg=1.11 M=.5516 Nbv=1.6989 N=1 Bv=8.1 Fc=.5 Ikf=0 Ibv=20.245m Is=880.5E-18 Xti=3) 
.model D1N750 D(Vj=.653 Cjo=175p Rs=.25 Eg=1.11 M=.5516 Nbv=1.6989 N=1 Bv=8.1 Fc=.5 Ikf=0 Ibv=20.245m Is=980.4E-18 Xti=3) 

* Dc analysis (varying Vin from -5 to 5 in steps of 0.01)
.ac dec 10 0.01 1Meg

* control statements
.control 
run
*white background set 
color0=white 
* black grid and text (only needed with X11, automatic with MS Win) 
set color1=yellow

* plotting waveforms
plot v(2) v(1)
*hardcopy xyPlot.ps v(1) v(2)
meas tran rptp pp v(2) from=10m to=40m
.endc


.end
