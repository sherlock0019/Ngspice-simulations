Full wave rectifier
*200030033_Q3a
V1 a 0 dc 0 Sin(0 2.5 1k 0 0 0)
D1 a b D1N750
D2 0 b D1N750
D3 c a D1N750
D4 c 0 D1N750
RL b c 1Meg
.model D1N750 D(Vj=.75 Cjo=175p Rs=.25 Eg=1.11 M=.5516 Nbv=1.6989 N=1 Bv=8.1 Fc=.5 Ikf=0 Ibv=20.245m Is=880.5E-18 Xti=3)
.tran 0.01ms 1ms

*control statements
.control
run

*white background
set color0=white
* black grid and text (only needed with X11, automatic with MS Win)
set color1=black
* wider grid and plot lines
set xbrushwidth=2

plot v(b,c) v(a)
.endc
.end

