Vin 2 1 Sin(0 16.9 50 0 0 0)
R1 1 4 0.01
vd1 4 5 0
vd2 3 6 0
.model 1N4001 D(Is=14.11n N=1.984 Rs=33.89m Ikf=94.81 Xti=3 Eg=1.11 Cjo=25.89p M=.44 Vj=.3245 Fc=.5 Bv=75 Ibv=10u Tt=5.7u Iave=1 Vpk=50 mfg=GI)

d1 5 3 1N4001
d2 2 3 1N4001
d3 0 2 1N4001
d4 0 5 1N4001
c1 6 0 3m
Rload 6 0 47
.tran 0.001s 0.1s 
.control 
 run 
*white background 
set color0=white 
* black grid and text (only needed with X11, automatic with MS Win) 
set color1=black 
* wider grid and plot lines 
set xbrushwidth=2 
* plotting input and output voltages 
plot v(1,2) v(6) i(vd1) i(vd2)
.endc 
.end
