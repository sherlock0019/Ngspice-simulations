BJT Common Emitter Amplifier Characteristics
vin 4 0 dc
vcc 7 0 12v

r1 7 4 31.33k
r2 4 0 10k
rc 7 5 5k
re 6 0 1.99k

*Dummy voltage sources to measure currents
vc 1 5 dc=0
vb 3 6 dc=0
ve 2 4 dc=0

Q1 1 2 3 Q2N2222A

.MODEL Q2N2222A NPN(IS=8.11E-14 BF=205 VAF=113 IKF=0.5 ISE=1.06E-11 + NE=2 BR=4 VAR=24 IKR=0.225 RB=1.37 RE=0.343 RC=0.137 CJE=2.95E-11 + TF=3.97E-10 CJC=1.52E-11 TR=8.5E-8 XTB=1.5)

.dc vin 0 12 12 

.control
run
print v(3), v(1,3), i(vc), i(vb), i(ve)
.endc
.end
