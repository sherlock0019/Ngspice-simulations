I/V characteristics of RED, GREEN and BLUE

V1 1 0 dc 0
R1 1 2 10k
R2 1 3 10k
R3 1 4 10k
D1 2 5 red
D2 3 6 green
D3 4 7 blue
V2 5 0 dc=0
V3 6 0 dc=0
V4 7 0 dc=0

.model red D(Vj=.75 Cjo=175p Rs=.25 Eg=3.2 M=.5516 Nbv=1.6989 N=2.4 Bv=1.7 Fc=.5 Ikf=0 Ibv=20.245m Is=880.5E-18 Xti=3)
.model green D(Is=1e-19 Rs=1.5 N=1.5 Cjo=50p Iave=30m Vpk=5)
.model blue D(IS=93.1P RS=42M N=7.47 BV=5 IBV=30U CJO=2.97P VJ=.75 M=.333 TT=4.32U)
.dc V1 0.001 10 0.001

.control
run
plot log(V2#branch) vs v(2,5), log(V3#branch) vs v(3,6), log(V4#branch) vs v(4,7)
.endc
.end
