Q-2 transient response of opamp model to confirm its working as an amplifier with Vfb offset
C1 0 3 10n IC=0v
R1 4 5 2k
R2 5 0 1k
E1 1 2 6 0 1
G1 0 3 2 0 0.01
E2 4 0 3 0 1
*Giving a step input
Vin 1 0 Pulse(0 1 0 0 10 10 10) 
Voff 5 6 0.1v 
.tran 0.004ms 4ms

.control
run
*plotting input and output voltages
plot v(1) v(4)
.endc
.end
