Amplifier

Vcc 3 0 12
Vin 4 0 1
Vdc 1 2 0
Vdb 5 8 0
Vde 6 9 0
*Cb 4 5 1u
*Ce 9 0 1u
*Cc 1 7 1u
Rc 3 1 5k
R1 3 5 33k
R2 5 0 10k
Re 9 0 2k
*Rl 7 0 1k
Q1 2 8 6 Q2N2222A

.MODEL Q2N2222A NPN(IS=8.11E-14 BF=205 VAF=113 IKF=0.5 ISE=1.06E-11
+ NE=2 BR=4 VAR=24 IKR=0.225 RB=1.37 RE=0.343 RC=0.137 CJE=2.95E-11
+ TF=3.97E-10 CJC=1.52E-11 TR=8.5E-8 XTB=1.5)

.control
op
dc vin 0 1 0.1
run

set color0=black
set color1=white
set xbrushwidth=2

plot i(Vdc)
plot i(Vdb)
plot i(Vde)
plot v(6)
plot v(1)
print i(8)
print i(6)
*plot v(7)
.endc
.end
